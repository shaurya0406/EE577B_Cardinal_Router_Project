`timescale 1ns/1ps
module cardinal_router (
  input  wire clk,
  input  wire reset
  // TODO: add channel I/O ports per spec
);
// TODO: RTL
endmodule
