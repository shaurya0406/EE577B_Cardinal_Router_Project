`timescale 1ns/1ps
module cardinal_nic (
  input  wire clk,
  input  wire reset
  // TODO: add processor & router-facing ports per spec
);
// TODO: RTL
endmodule
