`timescale 1ns/1ps
module router_tb;
  reg clk=0, reset=1;
  always #5 clk = ~clk;
  initial begin
    repeat (2) @(posedge clk);
    reset = 0;
    repeat (20) @(posedge clk);
    $finish;
  end
  cardinal_router dut(.clk(clk), .reset(reset));
endmodule
