`timescale 1ns/1ps
module cardinal_router_node (
  input  wire clk,
  input  wire reset
  // TODO: cw/ccw/pe ports
);
// TODO
endmodule
